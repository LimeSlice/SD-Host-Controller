module sd_receive (sd_clk, );


    wire [135:0] response;

    // multiple response types, either 48 bits or 136 bits


endmodule
